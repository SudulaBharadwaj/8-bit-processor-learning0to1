`timescale 1ns / 1ps


module NOT(
    input a,
    output op
    );
    assign op= ~a;
endmodule
